`timescale 1ns/1ps // Definir escala de tiempo
module ALU_TB();

// === Señales ===

//Registros
reg [31:0]xInput, yInput;
reg [4:0]sa_alu_tb;
reg [3:0]IN_OP;
//Conexiones
wire ZF_ALU_OUT;
wire [31:0]reOutput;
//Instancia
ALU alu(.sel(IN_OP),.zf(ZF_ALU_OUT),.x32bit(xInput[31:0]),.y32bit(yInput[31:0]),.shiftAmount(sa_alu_tb[4:0]),.res32bit(reOutput[31:0]));

// === Patrones de pruebas ===

initial
	begin
	IN_OP = 4'b0000; // Suma
	xInput[31:0] = 32'b00000000000000000000000011111111;
	yInput[31:0] = 32'b00000000000000000000000000000001;
	#10;
	
	xInput[31:0] = 32'b11111111111111111111111111111111;
	yInput[31:0] = 32'b11111111111111111111111111111111;
	#10;
	
	IN_OP = 4'b0001; // Resta
	
	xInput[31:0] = 32'b00000000000000000000000011111111;
	yInput[31:0] = 32'b00000000000000000000000000000001;
	#10;	
	
	xInput[31:0] = 32'b00000000000000000000000000000001;
	yInput[31:0] = 32'b11111111111111111111111111111111;
	#10;
	
	IN_OP = 4'b0010; // Multiplicacion
	
	xInput[31:0] = 32'b00000000000000000000000011111111;
	yInput[31:0] = 32'b00000000000000000000000000000001;
	#10;
	
	xInput[31:0] = 32'b00000000000000001111111111111111;
	yInput[31:0] = 32'b00000000000000001111111111111111;
	#10;

	IN_OP = 4'b0011; // Division
	
	xInput[31:0] = 32'b00000000000000000000000011111111;
	yInput[31:0] = 32'b00000000000000000000000000000001;
	#10;

	xInput[31:0] = 32'b00000000000000001111111111111111;
	yInput[31:0] = 32'b00000000000000000000000011111111;
	#10;

	IN_OP = 4'b0100; // AND
	
	xInput[31:0] = 32'b00000000000000000000000011111111;
	yInput[31:0] = 32'b00000000000000000000000000000001;
	#10;
	
	xInput[31:0] = 32'b11111111111111111111111111111111;
	yInput[31:0] = 32'b11111111111111111111111111111111;
	#10;
	
	IN_OP = 4'b0101; // OR
	
	xInput[31:0] = 32'b00000000000000000000000011111111;
	yInput[31:0] = 32'b00000000000000000000000000000001;
	#10;
	
	xInput[31:0] = 32'b11111111111111111111111111111111;
	yInput[31:0] = 32'b11111111111111111111111111111111;
	#10;
	
	IN_OP = 4'b0110; // NOR
	
	xInput[31:0] = 32'b00000000000000000000000011111111;
	yInput[31:0] = 32'b00000000000000000000000000000001;
	#10;
	
	xInput[31:0] = 32'b11111111111111111111111111111111;
	yInput[31:0] = 32'b11111111111111111111111111111111;
	#10;
	
	IN_OP = 4'b0111; // SLL
	
	sa_alu_tb[4:0] = 5'b00001; // left shift amount
	yInput[31:0] = 32'b00000000000000000000000000000001;
	#10;
	
	sa_alu_tb[4:0] = 5'b00001; // left shift amount
	yInput[31:0] = 32'b11111111111111111111111111111111;
	#10;
	
	IN_OP = 4'b1000; // SRL

	sa_alu_tb[4:0] = 5'b00001; // right shift amount
	yInput[31:0] = 32'b00000000000000000000000000000001;
	#10;

	sa_alu_tb[4:0] = 5'b00001; // right shift amount
	yInput[31:0] = 32'b11111111111111111111111111111111;
	#10;

	IN_OP = 4'b1001; // SLT
	
	xInput[31:0] = 32'b00000000000000000000000011111111;
	yInput[31:0] = 32'b00000000000000000000000000000001;
	#10;
	
	xInput[31:0] = 32'b11111111111111111111111111111111;
	yInput[31:0] = 32'b11111111111111111111111111111111;
	#10;
		
	IN_OP = 4'b1010; // XOR
	
	xInput[31:0] = 32'b00000000000000000000000011111111;
	yInput[31:0] = 32'b00000000000000000000000000000001;
	#10;
	
	xInput[31:0] = 32'b11111111111111111111111111111111;
	yInput[31:0] = 32'b11111111111111111111111111111111;
	#10;

	$stop;
	end
endmodule
